LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY EA IS	--Extensor Aritmético
	PORT (B: IN STD_LOGIC;
			S: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			SAIDA: OUT STD_LOGIC);
END;

ARCHITECTURE arch OF EA IS

SIGNAL aux: STD_LOGIC_VECTOR (2 DOWNTO 0);

BEGIN
	aux(0) <= S(3) AND B;
	aux(1) <= NOT S(2) AND NOT S(1) AND NOT S(0) AND B;
	aux(2) <= NOT S(3) AND NOT S(2) AND NOT S(1) AND S(0) AND NOT B;

	SAIDA <= aux(2) OR aux(1) OR aux(0);
END arch;